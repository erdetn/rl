// Copyright(C) 2022 Erdet Nasufi. All rights reserved.

module geometry

